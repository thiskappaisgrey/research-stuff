module test(
        input i_a,
        input i_b,
        output o_c
);
        
        assign o_c = i_a ^ i_b;
endmodule
